library ieee;
use ieee.std_logic_1164.all;

entity testbench is
end entity;

architecture bhv of testbench is

component AFG is
	port (Rx,clk, reset : in std_logic;
			outp : out std_logic_vector (7 downto 0));
end component AFG;
signal Rx, reset: std_logic:='1';
signal clk: std_logic:='0';
signal outp: std_logic_vector(7 downto 0);
begin
AFG1: AFG port map(Rx=>Rx, clk=>clk, reset=>reset, outp=>outp);

clk<= not clk after 20 ns;
reset<='0' after 10us;

pr:process
begin
rx<='1'; wait for 208 us;
rx <= '0'; wait for 104 us;--0
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--1
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--2
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--3
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--4
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--5
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--6
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--7
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--8
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--9
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--10
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--11
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--12
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--13
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--14
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--15
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--16
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--17
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--18
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--19
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--20
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--21
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--22
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--23
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;

rx <= '0'; wait for 104 us;--25
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--26
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '0'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
rx <= '0'; wait for 104 us;--27
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 936 us;
rx <= '0'; wait for 104 us;--24
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '0'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
        rx <= '1'; wait for 104 us;
		  rx <= '1'; wait for 1040 us;
end process;

end bhv;